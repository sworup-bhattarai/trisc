module two2one #(parameter N=4) 
  ( 
   input [N-1:0] A, B,   //declare data inputs 
   input S,   //declare select input 
   output [N-1:0] Y  //declare output 
  ); 
   assign Y = S==0 ? A : B; //select input 
  endmodule 